library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.STD_LOGIC_SIGNED.ALL;
use IEEE.NUMERIC_STD.ALL;

ENTITY ALU IS
	PORT(
	A1 : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
	A2 : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
	ALU_CONTROL : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
	ALU_RESULT : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
	ZERO : OUT STD_LOGIC;
	OVERFLOW : OUT STD_LOGIC
	);	
END ALU;

ARCHITECTURE Behavioral OF ALU IS
	SIGNAL RESULTX : STD_LOGIC_VECTOR(31 DOWNTO 0);
	SIGNAL RESULTP : STD_LOGIC_VECTOR(31 DOWNTO 0);
	SIGNAL C31_IN : std_logic;
	SIGNAL C31_OUT : std_logic;
BEGIN
	
	PROCESS(A1, A2, ALU_CONTROL)
	BEGIN
		CASE ALU_CONTROL IS
			WHEN "001" =>  -- ADDITION
				RESULTX <= STD_LOGIC_VECTOR(UNSIGNED(A1) + UNSIGNED(A2));
				RESULTP <= ("0" & A1(30 DOWNTO 0) + A2(30 DOWNTO 0));
				C31_IN <= RESULTP(31);
				C31_OUT <= ( (A1(31) XOR A2(31)) AND C31_IN) OR A1(31);
				OVERFLOW <= C31_IN XOR C31_OUT;
			WHEN "011" =>	-- SUB
				RESULTX <= STD_LOGIC_VECTOR(UNSIGNED(A1) - UNSIGNED(A2));
				RESULTP <= ("0" & A1(30 DOWNTO 0) + A2(30 DOWNTO 0));
				C31_IN <= RESULTP(31);
				C31_OUT <= ( (A1(31) XOR A2(31)) AND C31_IN) OR A1(31);
				OVERFLOW <= C31_IN XOR C31_OUT;
			WHEN "111" =>  -- AND
				RESULTX <= A1 AND A2;
				OVERFLOW <= '0';
			WHEN "010" =>  -- OR
				RESULTX <= A1 OR A2;
				OVERFLOW <= '0';
			WHEN OTHERS => 
			    RESULTX <= "00000000000000000000000000000000";
			    OVERFLOW <= '0';	   
		
		END CASE;
-- The reason i used a signal[RESULTX] to sore the output not dircetly store it in
-- "ALU_RESULT" because i will need to read it to decide the value of "ZERO"
-- and it's not possible to read an output
			
	END PROCESS;
	
	ALU_RESULT <= RESULTX;	   
	ZERO <= '1' WHEN RESULTX = "00000000000000000000000000000000" ELSE
		'0';

END Behavioral;
