LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.NUMERIC_STD.ALL;

ENTITY RegisterFile IS
	PORT(
	ReadRegister1 : IN STD_LOGIC_VECTOR (4 DOWNTO 0);
	ReadRegister2 : IN STD_LOGIC_VECTOR (4 DOWNTO 0);
	WriteRegister : IN STD_LOGIC_VECTOR (4 DOWNTO 0);
	RegWrite : IN STD_LOGIC;
	WriteData : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
	ReadData1 :	OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
	ReadData2 :	OUT STD_LOGIC_VECTOR (31 DOWNTO 0)
	);
END RegisterFile;

ARCHITECTURE Behavioral OF RegisterFile IS

	
	TYPE reg_file_type IS ARRAY(0 TO 31) OF
		STD_LOGIC_VECTOR(31 DOWNTO 0);
	
	
		
		
		
		
	SIGNAL array_reg : reg_file_type := ( 	"00000000000000000000000000000000",   --$zero 
											"00010001000100010001000100010001",   --$at
											"00100010001000100010001000100010",   --$v0
											"00110011001100110011001100110011",   --$v1
											"01000100010001000100010001000100",   --$a0
											"01010101010101010101010101010101",   --$a1
											"01100110011001100110011001100110",   --$a2
											"01110111011101110111011101110111",   --$a3
											"10001000100010001000100010001000",   --$t0
											"10011001100110011001100110011001",   --$t1
											"10101010101010101010101010101010",   --$t2
											"10111011101110111011101110111011",   --$t3
											"11001100110011001100110011001100",   --$t4
											"11011101110111011101110111011101",   --$t5
											"11101110111011101110111011101110",   --$t6
											"11111111111111111111111111111111",   --$t7
											"00000000000000000000000000000000",   --$s0
											"00010001000100010001000100010001",   --$s1
											"00100010001000100010001000100010",   --$s2
											"00110011001100110011001100110011",   --$s3
											"01000100010001000100010001000100",   --$s4
											"01010101010101010101010101010101",   --$s5
											"01100110011001100110011001100110",   --$s6
											"01110111011101110111011101110111",   --$s7
											"10001000100010001000100010001000",   --$t8
											"10011001100110011001100110011001",   --$t9
											"10101010101010101010101010101010",   --$k0
											"10111011101110111011101110111011",   --$k1
											"00010000000010000000000000000000",   --$gp
											"01101111111111111111000111101100",   --$sp
											"11101110111011101110111011101110",   --$fp
											"11111111111111111111111111111111"    --$ra
											);
BEGIN 
	PROCESS(RegWrite)
	BEGIN
		IF( RegWrite = '1' ) THEN
			array_reg(TO_INTEGER(UNSIGNED(WriteRegister))) <= WriteData;
		END IF;
	END PROCESS;  
				 -- i converted them to unsigned and to integer so i can use them as an index to the array
	ReadData1 <= array_reg(TO_INTEGER(UNSIGNED(ReadRegister1)));
	ReadData2 <= array_reg(TO_INTEGER(UNSIGNED(ReadRegister2)));
	
END Behavioral;
