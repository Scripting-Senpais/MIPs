library IEEE;
use IEEE.STD_LOGIC_1164.all;

entity MIPs is
	 port(
		 clk : in STD_LOGIC;
		 reset : in STD_LOGIC
	     );
end MIPs;

		 --just testing

architecture MIPs of MIPs is
begin



end MIPs;
